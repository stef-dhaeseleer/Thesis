`timescale 1ns / 1ps
`define RESET_TIME 25
`define CLK_PERIOD 10
`define CLK_HALF 5
`define EOF 32'hFFFF_FFFF 
`define NULL 0 

`include "des/des_pipelined.v"

// iverilog tb/tb_des_pipelined_automatic.v
// vvp a.out
// open -a gtkwave tb/vcd/tb_des_pipelined.vcd

module tb_des_pipelined();
    
    reg     clk;
    reg     rst_n;
    reg     start;
    reg [1:64] message;
    reg [1:768] round_keys;
    wire output_valid;
    wire [1:64] result;

    reg [1:64] expected;

    reg [14:0] nb_tests, nb_correct;
        
    //Instantiating montgomery module
    des_encryption_pipelined des_encryption_instance( 
            .clk            (clk         ),
            .rst_n          (rst_n       ),
            .start          (start       ),
            .message        (message     ),
            .round_keys     (round_keys  ),
            .output_valid   (output_valid),
            .result         (result      ));

    //Generate a clock
    initial begin
        clk = 0;
        forever #`CLK_HALF clk = ~clk;
    end
    
    //Reset
    initial begin
        rst_n = 0;
        #`RESET_TIME rst_n = 1;
    end
    
    //Test data
    initial begin

        $dumpfile("tb/vcd/tb_des_pipelined.vcd");
        $dumpvars(0, tb_des_pipelined);

        

        #`RESET_TIME

        // Init side parameters
        nb_tests <= 15'd0;
        nb_correct <= 15'd0;
                               
        #`CLK_PERIOD;

        // Wait until rising clock, read stimulus 
        @(posedge clk) 

            start<=1;
            #`CLK_PERIOD;
            start<=0;
            
            wait (output_valid==1);

            #`CLK_PERIOD;   // need this to check the result at the end of the done cycle and not at the start!

            nb_tests <= nb_tests + 1;
            nb_correct <= nb_correct + (expected - result == 64'h0);
                 
        $display("");
        $display("Correct tests: %d/%d", nb_correct, nb_tests);

        #`CLK_PERIOD;
        #`CLK_PERIOD;
  
        //r = $fcloser(file); 
        
        $finish;

    end
           
endmodule