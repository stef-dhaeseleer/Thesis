`timescale 1ns / 1ps
`define RESET_TIME 25
`define CLK_PERIOD 10
`define CLK_HALF 5
`define EOF 32'hFFFF_FFFF 
`define NULL 0 

`include "des/des_pipelined.v"

// iverilog tb/tb_des_pipelined_manual.v
// vvp a.out
// open -a gtkwave tb/vcd/tb_des_pipelined_manual.vcd

module tb_des_pipelined();
    
    reg     clk;
    reg     rst_n;
    reg     start;
    reg [1:64] message;
    reg [1:768] round_keys;
    wire output_valid;
    wire [1:64] result;

    reg [1:64] expected;

    reg [14:0] nb_tests, nb_correct;

    reg [1:64] message1;
    reg [1:64] expected1;
    reg [1:64] message2;
    reg [1:64] expected2;
    reg [1:64] message3;
    reg [1:64] expected3;
    reg [1:64] message4;
    reg [1:64] expected4;
    reg [1:64] message5;
    reg [1:64] expected5;
    reg [1:64] message6;
    reg [1:64] expected6;
    reg [1:64] message7;
    reg [1:64] expected7;
    reg [1:64] message8;
    reg [1:64] expected8;
    reg [1:64] message9;
    reg [1:64] expected9;
    reg [1:64] message10;
    reg [1:64] expected10;
    reg [1:64] message11;
    reg [1:64] expected11;
    reg [1:64] message12;
    reg [1:64] expected12;
    reg [1:64] message13;
    reg [1:64] expected13;
    reg [1:64] message14;
    reg [1:64] expected14;
    reg [1:64] message15;
    reg [1:64] expected15;
    reg [1:64] message16;
    reg [1:64] expected16;
    reg [1:64] message17;
    reg [1:64] expected17;
    reg [1:64] message18;
    reg [1:64] expected18;
    reg [1:64] message19;
    reg [1:64] expected19;
    reg [1:64] message20;
    reg [1:64] expected20;
    reg [1:64] message21;
    reg [1:64] expected21;
    reg [1:64] message22;
    reg [1:64] expected22;
    reg [1:64] message23;
    reg [1:64] expected23;
    reg [1:64] message24;
    reg [1:64] expected24;
    reg [1:64] message25;
    reg [1:64] expected25;
    reg [1:64] message26;
    reg [1:64] expected26;
    reg [1:64] message27;
    reg [1:64] expected27;
    reg [1:64] message28;
    reg [1:64] expected28;
    reg [1:64] message29;
    reg [1:64] expected29;
    reg [1:64] message30;
    reg [1:64] expected30;
    reg [1:64] message31;
    reg [1:64] expected31;
    reg [1:64] message32;
    reg [1:64] expected32;
    reg [1:64] message33;
    reg [1:64] expected33;
    reg [1:64] message34;
    reg [1:64] expected34;
    reg [1:64] message35;
    reg [1:64] expected35;
    reg [1:64] message36;
    reg [1:64] expected36;
    reg [1:64] message37;
    reg [1:64] expected37;
    reg [1:64] message38;
    reg [1:64] expected38;
    reg [1:64] message39;
    reg [1:64] expected39;
    reg [1:64] message40;
    reg [1:64] expected40;
    reg [1:64] message41;
    reg [1:64] expected41;
    reg [1:64] message42;
    reg [1:64] expected42;
    reg [1:64] message43;
    reg [1:64] expected43;
    reg [1:64] message44;
    reg [1:64] expected44;
    reg [1:64] message45;
    reg [1:64] expected45;
    reg [1:64] message46;
    reg [1:64] expected46;
    reg [1:64] message47;
    reg [1:64] expected47;
    reg [1:64] message48;
    reg [1:64] expected48;
    reg [1:64] message49;
    reg [1:64] expected49;
    reg [1:64] message50;
    reg [1:64] expected50;
    reg [1:64] message51;
    reg [1:64] expected51;
    reg [1:64] message52;
    reg [1:64] expected52;
    reg [1:64] message53;
    reg [1:64] expected53;
    reg [1:64] message54;
    reg [1:64] expected54;
    reg [1:64] message55;
    reg [1:64] expected55;
    reg [1:64] message56;
    reg [1:64] expected56;
    reg [1:64] message57;
    reg [1:64] expected57;
    reg [1:64] message58;
    reg [1:64] expected58;
    reg [1:64] message59;
    reg [1:64] expected59;
    reg [1:64] message60;
    reg [1:64] expected60;
    reg [1:64] message61;
    reg [1:64] expected61;
    reg [1:64] message62;
    reg [1:64] expected62;
    reg [1:64] message63;
    reg [1:64] expected63;
    reg [1:64] message64;
    reg [1:64] expected64;
    reg [1:64] message65;
    reg [1:64] expected65;
    reg [1:64] message66;
    reg [1:64] expected66;
    reg [1:64] message67;
    reg [1:64] expected67;
    reg [1:64] message68;
    reg [1:64] expected68;
    reg [1:64] message69;
    reg [1:64] expected69;
    reg [1:64] message70;
    reg [1:64] expected70;
    reg [1:64] message71;
    reg [1:64] expected71;
    reg [1:64] message72;
    reg [1:64] expected72;
    reg [1:64] message73;
    reg [1:64] expected73;
    reg [1:64] message74;
    reg [1:64] expected74;
    reg [1:64] message75;
    reg [1:64] expected75;
    reg [1:64] message76;
    reg [1:64] expected76;
    reg [1:64] message77;
    reg [1:64] expected77;
    reg [1:64] message78;
    reg [1:64] expected78;
    reg [1:64] message79;
    reg [1:64] expected79;
    reg [1:64] message80;
    reg [1:64] expected80;
    reg [1:64] message81;
    reg [1:64] expected81;
    reg [1:64] message82;
    reg [1:64] expected82;
    reg [1:64] message83;
    reg [1:64] expected83;
    reg [1:64] message84;
    reg [1:64] expected84;
    reg [1:64] message85;
    reg [1:64] expected85;
    reg [1:64] message86;
    reg [1:64] expected86;
    reg [1:64] message87;
    reg [1:64] expected87;
    reg [1:64] message88;
    reg [1:64] expected88;
    reg [1:64] message89;
    reg [1:64] expected89;
    reg [1:64] message90;
    reg [1:64] expected90;
    reg [1:64] message91;
    reg [1:64] expected91;
    reg [1:64] message92;
    reg [1:64] expected92;
    reg [1:64] message93;
    reg [1:64] expected93;
    reg [1:64] message94;
    reg [1:64] expected94;
    reg [1:64] message95;
    reg [1:64] expected95;
    reg [1:64] message96;
    reg [1:64] expected96;
    reg [1:64] message97;
    reg [1:64] expected97;
    reg [1:64] message98;
    reg [1:64] expected98;
    reg [1:64] message99;
    reg [1:64] expected99;
    reg [1:64] message100;
    reg [1:64] expected100;
    reg [1:64] message101;
    reg [1:64] expected101;
    reg [1:64] message102;
    reg [1:64] expected102;
    reg [1:64] message103;
    reg [1:64] expected103;
    reg [1:64] message104;
    reg [1:64] expected104;
    reg [1:64] message105;
    reg [1:64] expected105;
    reg [1:64] message106;
    reg [1:64] expected106;
    reg [1:64] message107;
    reg [1:64] expected107;
    reg [1:64] message108;
    reg [1:64] expected108;
    reg [1:64] message109;
    reg [1:64] expected109;
    reg [1:64] message110;
    reg [1:64] expected110;
    reg [1:64] message111;
    reg [1:64] expected111;
    reg [1:64] message112;
    reg [1:64] expected112;
    reg [1:64] message113;
    reg [1:64] expected113;
    reg [1:64] message114;
    reg [1:64] expected114;
    reg [1:64] message115;
    reg [1:64] expected115;
    reg [1:64] message116;
    reg [1:64] expected116;
    reg [1:64] message117;
    reg [1:64] expected117;
    reg [1:64] message118;
    reg [1:64] expected118;
    reg [1:64] message119;
    reg [1:64] expected119;
    reg [1:64] message120;
    reg [1:64] expected120;
    reg [1:64] message121;
    reg [1:64] expected121;
    reg [1:64] message122;
    reg [1:64] expected122;
    reg [1:64] message123;
    reg [1:64] expected123;
    reg [1:64] message124;
    reg [1:64] expected124;
    reg [1:64] message125;
    reg [1:64] expected125;
    reg [1:64] message126;
    reg [1:64] expected126;
    reg [1:64] message127;
    reg [1:64] expected127;
    reg [1:64] message128;
    reg [1:64] expected128;
        
    //Instantiating montgomery module
    des_encryption_pipelined des_encryption_instance( 
            .clk            (clk         ),
            .rst_n          (rst_n       ),
            .start          (start       ),
            .message        (message     ),
            .round_keys     (round_keys  ),
            .output_valid   (output_valid),
            .result         (result      ));

    //Generate a clock
    initial begin
        clk = 0;
        forever #`CLK_HALF clk = ~clk;
    end
    
    //Reset
    initial begin
        rst_n = 0;
        #`RESET_TIME rst_n = 1;
    end
    
    //Test data
    initial begin

        $dumpfile("tb/vcd/tb_des_pipelined_manual.vcd");
        $dumpvars(0, tb_des_pipelined);

        #`RESET_TIME
    
        round_keys <= 768'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        
        message1 <= 64'b1001010111111000101001011110010111011101001100011101100100000000;
        expected1 <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
        message2 <= 64'b1101110101111111000100100001110010100101000000010101011000011001;
        expected2 <= 64'b0100000000000000000000000000000000000000000000000000000000000000;
        message3 <= 64'b0010111010000110010100110001000001001111001110000011010011101010;
        expected3 <= 64'b0010000000000000000000000000000000000000000000000000000000000000;
        message4 <= 64'b0100101111010011100010001111111101101100110110000001110101001111;
        expected4 <= 64'b0001000000000000000000000000000000000000000000000000000000000000;
        message5 <= 64'b0010000010111001111001110110011110110010111110110001010001010110;
        expected5 <= 64'b0000100000000000000000000000000000000000000000000000000000000000;
        message6 <= 64'b0101010101010111100100111000000011010111011100010011100011101111;
        expected6 <= 64'b0000010000000000000000000000000000000000000000000000000000000000;
        message7 <= 64'b0110110011000101110111101111101010101111000001000101000100101111;
        expected7 <= 64'b0000001000000000000000000000000000000000000000000000000000000000;
        message8 <= 64'b0000110110011111001001111001101110100101110110000111001001100000;
        expected8 <= 64'b0000000100000000000000000000000000000000000000000000000000000000;
        message9 <= 64'b1101100100000011000110110000001001110001101111010101101000001010;
        expected9 <= 64'b0000000010000000000000000000000000000000000000000000000000000000;
        message10 <= 64'b0100001001000010010100001011001101111100001111011101100101010001;
        expected10 <= 64'b0000000001000000000000000000000000000000000000000000000000000000;
        message11 <= 64'b1011100000000110000110110111111011001101100110100010000111100101;
        expected11 <= 64'b0000000000100000000000000000000000000000000000000000000000000000;
        message12 <= 64'b1111000101011101000011110010100001101011011001011011110100101000;
        expected12 <= 64'b0000000000010000000000000000000000000000000000000000000000000000;
        message13 <= 64'b1010110111010000110011001000110101101110010111011110101110100001;
        expected13 <= 64'b0000000000001000000000000000000000000000000000000000000000000000;
        message14 <= 64'b1110011011010101111110000010011101010010101011010110001111010001;
        expected14 <= 64'b0000000000000100000000000000000000000000000000000000000000000000;
        message15 <= 64'b1110110010111111111000111011110100111111010110010001101001011110;
        expected15 <= 64'b0000000000000010000000000000000000000000000000000000000000000000;
        message16 <= 64'b1111001101010110100000110100001101111001110100010110010111001101;
        expected16 <= 64'b0000000000000001000000000000000000000000000000000000000000000000;
        message17 <= 64'b0010101110011111100110000010111100100000000000110111111110101001;
        expected17 <= 64'b0000000000000000100000000000000000000000000000000000000000000000;
        message18 <= 64'b1000100010011101111000000110100010100001011011110000101111100110;
        expected18 <= 64'b0000000000000000010000000000000000000000000000000000000000000000;
        message19 <= 64'b1110000110011110001001110101110110000100011010100001001010011000;
        expected19 <= 64'b0000000000000000001000000000000000000000000000000000000000000000;
        message20 <= 64'b0011001010011010100011101101010100100011110101110001101011101100;
        expected20 <= 64'b0000000000000000000100000000000000000000000000000000000000000000;
        message21 <= 64'b1110011111111100111000100010010101010111110100100011110010010111;
        expected21 <= 64'b0000000000000000000010000000000000000000000000000000000000000000;
        message22 <= 64'b0001001010101001111101011000000101111111111100101101011001011101;
        expected22 <= 64'b0000000000000000000001000000000000000000000000000000000000000000;
        message23 <= 64'b1010010010000100110000111010110100111000110111001001110000011001;
        expected23 <= 64'b0000000000000000000000100000000000000000000000000000000000000000;
        message24 <= 64'b1111101111100000000010101000101000011110111110001010110101110010;
        expected24 <= 64'b0000000000000000000000010000000000000000000000000000000000000000;
        message25 <= 64'b0111010100001101000001111001010000000111010100100001001101100011;
        expected25 <= 64'b0000000000000000000000001000000000000000000000000000000000000000;
        message26 <= 64'b0110010011111110111011011001110001110010010011000010111110101111;
        expected26 <= 64'b0000000000000000000000000100000000000000000000000000000000000000;
        message27 <= 64'b1111000000101011001001100011101100110010100011100010101101100000;
        expected27 <= 64'b0000000000000000000000000010000000000000000000000000000000000000;
        message28 <= 64'b1001110101100100010101010101101010011010000100001011100001010010;
        expected28 <= 64'b0000000000000000000000000001000000000000000000000000000000000000;
        message29 <= 64'b1101000100000110111111110000101111101101010100100101010111010111;
        expected29 <= 64'b0000000000000000000000000000100000000000000000000000000000000000;
        message30 <= 64'b1110000101100101001011000110101100010011100011000110010010100101;
        expected30 <= 64'b0000000000000000000000000000010000000000000000000000000000000000;
        message31 <= 64'b1110010000101000010110000001000110000110111011001000111101000110;
        expected31 <= 64'b0000000000000000000000000000001000000000000000000000000000000000;
        message32 <= 64'b1010111010110101111101011110110111100010001011010001101000110110;
        expected32 <= 64'b0000000000000000000000000000000100000000000000000000000000000000;
        message33 <= 64'b1110100101000011110101110101011010001010111011000000110001011100;
        expected33 <= 64'b0000000000000000000000000000000010000000000000000000000000000000;
        message34 <= 64'b1101111110011000110010000010011101101111010101001011000001001011;
        expected34 <= 64'b0000000000000000000000000000000001000000000000000000000000000000;
        message35 <= 64'b1011000101100000111001000110100000001111011011000110100101101111;
        expected35 <= 64'b0000000000000000000000000000000000100000000000000000000000000000;
        message36 <= 64'b1111101000000111010100101011000001111101100111000100101010111000;
        expected36 <= 64'b0000000000000000000000000000000000010000000000000000000000000000;
        message37 <= 64'b1100101000111010001010110000001101101101101111001000010100000010;
        expected37 <= 64'b0000000000000000000000000000000000001000000000000000000000000000;
        message38 <= 64'b0101111000001001000001010101000101111011101101011001101111001111;
        expected38 <= 64'b0000000000000000000000000000000000000100000000000000000000000000;
        message39 <= 64'b1000000101001110111010110011101110010001110110010000011100100110;
        expected39 <= 64'b0000000000000000000000000000000000000010000000000000000000000000;
        message40 <= 64'b0100110101001001110110110001010100110010100100011001110010011111;
        expected40 <= 64'b0000000000000000000000000000000000000001000000000000000000000000;
        message41 <= 64'b0010010111101011010111111100001111111000110011110000011000100001;
        expected41 <= 64'b0000000000000000000000000000000000000000100000000000000000000000;
        message42 <= 64'b1010101101101010001000001100000001100010000011010001110001101111;
        expected42 <= 64'b0000000000000000000000000000000000000000010000000000000000000000;
        message43 <= 64'b0111100111101001000011011011110010011000111110010010110011001010;
        expected43 <= 64'b0000000000000000000000000000000000000000001000000000000000000000;
        message44 <= 64'b1000011001101110110011101101110110000000011100101011101100001110;
        expected44 <= 64'b0000000000000000000000000000000000000000000100000000000000000000;
        message45 <= 64'b1000101101010100010100110110111100101111001111100110010010101000;
        expected45 <= 64'b0000000000000000000000000000000000000000000010000000000000000000;
        message46 <= 64'b1110101001010001110100111001011101010101100101011011100001101011;
        expected46 <= 64'b0000000000000000000000000000000000000000000001000000000000000000;
        message47 <= 64'b1100101011111111110001101010110001000101010000101101111000110001;
        expected47 <= 64'b0000000000000000000000000000000000000000000000100000000000000000;
        message48 <= 64'b1000110111010100010110100010110111011111100100000111100101101100;
        expected48 <= 64'b0000000000000000000000000000000000000000000000010000000000000000;
        message49 <= 64'b0001000000101001110101010101111010001000000011101100001011010000;
        expected49 <= 64'b0000000000000000000000000000000000000000000000001000000000000000;
        message50 <= 64'b0101110110000110110010110010001101100011100111011011111010101001;
        expected50 <= 64'b0000000000000000000000000000000000000000000000000100000000000000;
        message51 <= 64'b0001110100011100101010000101001110101110011111000000110001011111;
        expected51 <= 64'b0000000000000000000000000000000000000000000000000010000000000000;
        message52 <= 64'b1100111000110011001000110010100100100100100011110011001000101000;
        expected52 <= 64'b0000000000000000000000000000000000000000000000000001000000000000;
        message53 <= 64'b1000010000000101110100011010101111100010010011111011100101000010;
        expected53 <= 64'b0000000000000000000000000000000000000000000000000000100000000000;
        message54 <= 64'b1110011001000011110101111000000010010000110010100100001000000111;
        expected54 <= 64'b0000000000000000000000000000000000000000000000000000010000000000;
        message55 <= 64'b0100100000100010000110111001100100110111011101001000101000100011;
        expected55 <= 64'b0000000000000000000000000000000000000000000000000000001000000000;
        message56 <= 64'b1101110101111100000010111011110101100001111110101111110101010100;
        expected56 <= 64'b0000000000000000000000000000000000000000000000000000000100000000;
        message57 <= 64'b0010111110111100001010010001101001010111000011011011010111000100;
        expected57 <= 64'b0000000000000000000000000000000000000000000000000000000010000000;
        message58 <= 64'b1110000001111100001100001101011111100100111000100110111000010010;
        expected58 <= 64'b0000000000000000000000000000000000000000000000000000000001000000;
        message59 <= 64'b0000100101010011111000100010010110001110100011101001000010100001;
        expected59 <= 64'b0000000000000000000000000000000000000000000000000000000000100000;
        message60 <= 64'b0101101101110001000110111100010011001110111010111111001011101110;
        expected60 <= 64'b0000000000000000000000000000000000000000000000000000000000010000;
        message61 <= 64'b1100110000001000001111110001111001101101100111101000010111110110;
        expected61 <= 64'b0000000000000000000000000000000000000000000000000000000000001000;
        message62 <= 64'b1101001011111101100010000110011111010101000011010010110111111110;
        expected62 <= 64'b0000000000000000000000000000000000000000000000000000000000000100;
        message63 <= 64'b0000011011100111111010100010001011001110100100100111000010001111;
        expected63 <= 64'b0000000000000000000000000000000000000000000000000000000000000010;
        message64 <= 64'b0001011001101011010000001011010001001010101110100100101111010110;
        expected64 <= 64'b0000000000000000000000000000000000000000000000000000000000000001;
        message65 <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
        expected65 <= 64'b1001010111111000101001011110010111011101001100011101100100000000;
        message66 <= 64'b0100000000000000000000000000000000000000000000000000000000000000;
        expected66 <= 64'b1101110101111111000100100001110010100101000000010101011000011001;
        message67 <= 64'b0010000000000000000000000000000000000000000000000000000000000000;
        expected67 <= 64'b0010111010000110010100110001000001001111001110000011010011101010;
        message68 <= 64'b0001000000000000000000000000000000000000000000000000000000000000;
        expected68 <= 64'b0100101111010011100010001111111101101100110110000001110101001111;
        message69 <= 64'b0000100000000000000000000000000000000000000000000000000000000000;
        expected69 <= 64'b0010000010111001111001110110011110110010111110110001010001010110;
        message70 <= 64'b0000010000000000000000000000000000000000000000000000000000000000;
        expected70 <= 64'b0101010101010111100100111000000011010111011100010011100011101111;
        message71 <= 64'b0000001000000000000000000000000000000000000000000000000000000000;
        expected71 <= 64'b0110110011000101110111101111101010101111000001000101000100101111;
        message72 <= 64'b0000000100000000000000000000000000000000000000000000000000000000;
        expected72 <= 64'b0000110110011111001001111001101110100101110110000111001001100000;
        message73 <= 64'b0000000010000000000000000000000000000000000000000000000000000000;
        expected73 <= 64'b1101100100000011000110110000001001110001101111010101101000001010;
        message74 <= 64'b0000000001000000000000000000000000000000000000000000000000000000;
        expected74 <= 64'b0100001001000010010100001011001101111100001111011101100101010001;
        message75 <= 64'b0000000000100000000000000000000000000000000000000000000000000000;
        expected75 <= 64'b1011100000000110000110110111111011001101100110100010000111100101;
        message76 <= 64'b0000000000010000000000000000000000000000000000000000000000000000;
        expected76 <= 64'b1111000101011101000011110010100001101011011001011011110100101000;
        message77 <= 64'b0000000000001000000000000000000000000000000000000000000000000000;
        expected77 <= 64'b1010110111010000110011001000110101101110010111011110101110100001;
        message78 <= 64'b0000000000000100000000000000000000000000000000000000000000000000;
        expected78 <= 64'b1110011011010101111110000010011101010010101011010110001111010001;
        message79 <= 64'b0000000000000010000000000000000000000000000000000000000000000000;
        expected79 <= 64'b1110110010111111111000111011110100111111010110010001101001011110;
        message80 <= 64'b0000000000000001000000000000000000000000000000000000000000000000;
        expected80 <= 64'b1111001101010110100000110100001101111001110100010110010111001101;
        message81 <= 64'b0000000000000000100000000000000000000000000000000000000000000000;
        expected81 <= 64'b0010101110011111100110000010111100100000000000110111111110101001;
        message82 <= 64'b0000000000000000010000000000000000000000000000000000000000000000;
        expected82 <= 64'b1000100010011101111000000110100010100001011011110000101111100110;
        message83 <= 64'b0000000000000000001000000000000000000000000000000000000000000000;
        expected83 <= 64'b1110000110011110001001110101110110000100011010100001001010011000;
        message84 <= 64'b0000000000000000000100000000000000000000000000000000000000000000;
        expected84 <= 64'b0011001010011010100011101101010100100011110101110001101011101100;
        message85 <= 64'b0000000000000000000010000000000000000000000000000000000000000000;
        expected85 <= 64'b1110011111111100111000100010010101010111110100100011110010010111;
        message86 <= 64'b0000000000000000000001000000000000000000000000000000000000000000;
        expected86 <= 64'b0001001010101001111101011000000101111111111100101101011001011101;
        message87 <= 64'b0000000000000000000000100000000000000000000000000000000000000000;
        expected87 <= 64'b1010010010000100110000111010110100111000110111001001110000011001;
        message88 <= 64'b0000000000000000000000010000000000000000000000000000000000000000;
        expected88 <= 64'b1111101111100000000010101000101000011110111110001010110101110010;
        message89 <= 64'b0000000000000000000000001000000000000000000000000000000000000000;
        expected89 <= 64'b0111010100001101000001111001010000000111010100100001001101100011;
        message90 <= 64'b0000000000000000000000000100000000000000000000000000000000000000;
        expected90 <= 64'b0110010011111110111011011001110001110010010011000010111110101111;
        message91 <= 64'b0000000000000000000000000010000000000000000000000000000000000000;
        expected91 <= 64'b1111000000101011001001100011101100110010100011100010101101100000;
        message92 <= 64'b0000000000000000000000000001000000000000000000000000000000000000;
        expected92 <= 64'b1001110101100100010101010101101010011010000100001011100001010010;
        message93 <= 64'b0000000000000000000000000000100000000000000000000000000000000000;
        expected93 <= 64'b1101000100000110111111110000101111101101010100100101010111010111;
        message94 <= 64'b0000000000000000000000000000010000000000000000000000000000000000;
        expected94 <= 64'b1110000101100101001011000110101100010011100011000110010010100101;
        message95 <= 64'b0000000000000000000000000000001000000000000000000000000000000000;
        expected95 <= 64'b1110010000101000010110000001000110000110111011001000111101000110;
        message96 <= 64'b0000000000000000000000000000000100000000000000000000000000000000;
        expected96 <= 64'b1010111010110101111101011110110111100010001011010001101000110110;
        message97 <= 64'b0000000000000000000000000000000010000000000000000000000000000000;
        expected97 <= 64'b1110100101000011110101110101011010001010111011000000110001011100;
        message98 <= 64'b0000000000000000000000000000000001000000000000000000000000000000;
        expected98 <= 64'b1101111110011000110010000010011101101111010101001011000001001011;
        message99 <= 64'b0000000000000000000000000000000000100000000000000000000000000000;
        expected99 <= 64'b1011000101100000111001000110100000001111011011000110100101101111;
        message100 <= 64'b0000000000000000000000000000000000010000000000000000000000000000;
        expected100 <= 64'b1111101000000111010100101011000001111101100111000100101010111000;
        message101 <= 64'b0000000000000000000000000000000000001000000000000000000000000000;
        expected101 <= 64'b1100101000111010001010110000001101101101101111001000010100000010;
        message102 <= 64'b0000000000000000000000000000000000000100000000000000000000000000;
        expected102 <= 64'b0101111000001001000001010101000101111011101101011001101111001111;
        message103 <= 64'b0000000000000000000000000000000000000010000000000000000000000000;
        expected103 <= 64'b1000000101001110111010110011101110010001110110010000011100100110;
        message104 <= 64'b0000000000000000000000000000000000000001000000000000000000000000;
        expected104 <= 64'b0100110101001001110110110001010100110010100100011001110010011111;
        message105 <= 64'b0000000000000000000000000000000000000000100000000000000000000000;
        expected105 <= 64'b0010010111101011010111111100001111111000110011110000011000100001;
        message106 <= 64'b0000000000000000000000000000000000000000010000000000000000000000;
        expected106 <= 64'b1010101101101010001000001100000001100010000011010001110001101111;
        message107 <= 64'b0000000000000000000000000000000000000000001000000000000000000000;
        expected107 <= 64'b0111100111101001000011011011110010011000111110010010110011001010;
        message108 <= 64'b0000000000000000000000000000000000000000000100000000000000000000;
        expected108 <= 64'b1000011001101110110011101101110110000000011100101011101100001110;
        message109 <= 64'b0000000000000000000000000000000000000000000010000000000000000000;
        expected109 <= 64'b1000101101010100010100110110111100101111001111100110010010101000;
        message110 <= 64'b0000000000000000000000000000000000000000000001000000000000000000;
        expected110 <= 64'b1110101001010001110100111001011101010101100101011011100001101011;
        message111 <= 64'b0000000000000000000000000000000000000000000000100000000000000000;
        expected111 <= 64'b1100101011111111110001101010110001000101010000101101111000110001;
        message112 <= 64'b0000000000000000000000000000000000000000000000010000000000000000;
        expected112 <= 64'b1000110111010100010110100010110111011111100100000111100101101100;
        message113 <= 64'b0000000000000000000000000000000000000000000000001000000000000000;
        expected113 <= 64'b0001000000101001110101010101111010001000000011101100001011010000;
        message114 <= 64'b0000000000000000000000000000000000000000000000000100000000000000;
        expected114 <= 64'b0101110110000110110010110010001101100011100111011011111010101001;
        message115 <= 64'b0000000000000000000000000000000000000000000000000010000000000000;
        expected115 <= 64'b0001110100011100101010000101001110101110011111000000110001011111;
        message116 <= 64'b0000000000000000000000000000000000000000000000000001000000000000;
        expected116 <= 64'b1100111000110011001000110010100100100100100011110011001000101000;
        message117 <= 64'b0000000000000000000000000000000000000000000000000000100000000000;
        expected117 <= 64'b1000010000000101110100011010101111100010010011111011100101000010;
        message118 <= 64'b0000000000000000000000000000000000000000000000000000010000000000;
        expected118 <= 64'b1110011001000011110101111000000010010000110010100100001000000111;
        message119 <= 64'b0000000000000000000000000000000000000000000000000000001000000000;
        expected119 <= 64'b0100100000100010000110111001100100110111011101001000101000100011;
        message120 <= 64'b0000000000000000000000000000000000000000000000000000000100000000;
        expected120 <= 64'b1101110101111100000010111011110101100001111110101111110101010100;
        message121 <= 64'b0000000000000000000000000000000000000000000000000000000010000000;
        expected121 <= 64'b0010111110111100001010010001101001010111000011011011010111000100;
        message122 <= 64'b0000000000000000000000000000000000000000000000000000000001000000;
        expected122 <= 64'b1110000001111100001100001101011111100100111000100110111000010010;
        message123 <= 64'b0000000000000000000000000000000000000000000000000000000000100000;
        expected123 <= 64'b0000100101010011111000100010010110001110100011101001000010100001;
        message124 <= 64'b0000000000000000000000000000000000000000000000000000000000010000;
        expected124 <= 64'b0101101101110001000110111100010011001110111010111111001011101110;
        message125 <= 64'b0000000000000000000000000000000000000000000000000000000000001000;
        expected125 <= 64'b1100110000001000001111110001111001101101100111101000010111110110;
        message126 <= 64'b0000000000000000000000000000000000000000000000000000000000000100;
        expected126 <= 64'b1101001011111101100010000110011111010101000011010010110111111110;
        message127 <= 64'b0000000000000000000000000000000000000000000000000000000000000010;
        expected127 <= 64'b0000011011100111111010100010001011001110100100100111000010001111;
        message128 <= 64'b0000000000000000000000000000000000000000000000000000000000000001;
        expected128 <= 64'b0001011001101011010000001011010001001010101110100100101111010110;

        // Init side parameters
        nb_tests <= 15'd0;
        nb_correct <= 15'd0;
                               
        #`CLK_PERIOD;

        // Wait until rising clock, read stimulus 
        start<=1;
        message <= message1;
        #`CLK_PERIOD;
        //start<=0;
        message <= message2;
        #`CLK_PERIOD;
        message <= message3;
        #`CLK_PERIOD;
        message <= message4;
        #`CLK_PERIOD;
        message <= message5;
        #`CLK_PERIOD;
        message <= message6;
        #`CLK_PERIOD;
        message <= message7;
        #`CLK_PERIOD;
        message <= message8;
        #`CLK_PERIOD;
        message <= message9;
        #`CLK_PERIOD;
        message <= message10;
        #`CLK_PERIOD;
        message <= message11;
        #`CLK_PERIOD;
        message <= message12;
        #`CLK_PERIOD;
        message <= message13;
        #`CLK_PERIOD;
        message <= message14;
        #`CLK_PERIOD;
        message <= message15;
        #`CLK_PERIOD;
        message <= message16;
        #`CLK_PERIOD;
        message <= message17;
        #`CLK_PERIOD;
        message <= message18;
        #`CLK_PERIOD;

        message <= message19;
        #`CLK_PERIOD;

        message <= message20;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected1 - result == 64'h0);
        #`CLK_PERIOD;
        
        message <= message21;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected2 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message22;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected3 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message23;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected4 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message24;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected5 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message25;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected6 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message26;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected7 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message27;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected8 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message28;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected9 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message29;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected10 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message30;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected11 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message31;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected12 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message32;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected13 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message33;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected14 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message34;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected15 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message35;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected16 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message36;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected17 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message37;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected18 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message38;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected19 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message39;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected20 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message40;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected21 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message41;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected22 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message42;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected23 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message43;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected24 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message44;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected25 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message45;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected26 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message46;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected27 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message47;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected28 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message48;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected29 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message49;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected30 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message50;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected31 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message51;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected32 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message52;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected33 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message53;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected34 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message54;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected35 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message55;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected36 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message56;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected37 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message57;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected38 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message58;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected39 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message59;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected40 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message60;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected41 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message61;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected42 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message62;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected43 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message63;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected44 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message64;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected45 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message65;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected46 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message66;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected47 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message67;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected48 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message68;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected49 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message69;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected50 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message70;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected51 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message71;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected52 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message72;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected53 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message73;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected54 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message74;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected55 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message75;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected56 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message76;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected57 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message77;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected58 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message78;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected59 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message79;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected60 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message80;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected61 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message81;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected62 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message82;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected63 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message83;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected64 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message84;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected65 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message85;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected66 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message86;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected67 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message87;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected68 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message88;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected69 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message89;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected70 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message90;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected71 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message91;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected72 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message92;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected73 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message93;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected74 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message94;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected75 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message95;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected76 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message96;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected77 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message97;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected78 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message98;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected79 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message99;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected80 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message100;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected81 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message101;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected82 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message102;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected83 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message103;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected84 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message104;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected85 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message105;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected86 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message106;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected87 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message107;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected88 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message108;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected89 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message109;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected90 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message110;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected91 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message111;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected92 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message112;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected93 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message113;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected94 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message114;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected95 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message115;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected96 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message116;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected97 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message117;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected98 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message118;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected99 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message119;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected100 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message120;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected101 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message121;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected102 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message122;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected103 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message123;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected104 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message124;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected105 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message125;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected106 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message126;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected107 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message127;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected108 - result == 64'h0);
        #`CLK_PERIOD;

        message <= message128;
        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected109 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected110 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected111 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected112 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected113 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected114 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected115 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected116 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected117 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected118 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected119 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected120 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected121 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected122 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected123 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected124 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected125 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected126 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected127 - result == 64'h0);
        #`CLK_PERIOD;

        nb_tests <= nb_tests + 1;
        nb_correct <= nb_correct + (expected128 - result == 64'h0);
        #`CLK_PERIOD;

        $display("");
        $display("Correct tests: %d/%d", nb_correct, nb_tests);

        #`CLK_PERIOD;
        #`CLK_PERIOD;

    
        $finish;

    end
           
endmodule